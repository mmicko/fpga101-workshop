module led (
    output LED_B
);
    assign LED_B = 1'b0;
endmodule
